** Profile: "SCHEMATIC1-DC"  [ E:\PCB_ESP_CON_USB\Datasheets\INA157U\INA157_PSPICE_AIO\ina157-pspicefiles\schematic1\dc.sim ] 

** Creating circuit file "DC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../INA157.lib" 
* From [PSPICE NETLIST] section of F:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_VIN -20 20 0.01 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
